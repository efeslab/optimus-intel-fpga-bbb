`define MPF_CONF_SORT_READ_RESPONSES            1
`define MPF_CONF_PRESERVE_WRITE_MDATA           0
`define MPF_CONF_ENABLE_VC_MAP                  0
`define MPF_CONF_ENABLE_DYNAMIC_VC_MAPPING      0
`define MPF_CONF_ENABLE_LATENCY_QOS             0
`define MPF_CONF_ENFORCE_WR_ORDER               0
`define MPF_CONF_ENABLE_PARTIAL_WRITES          0
`define MPF_CONF_MERGE_DUPLICATE_READS          0
