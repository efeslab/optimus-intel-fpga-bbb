// RO
